`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/01/2023 03:48:05 PM
// Design Name: 
// Module Name: controlNode
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module controlNode(input logic clk, read_i, write_i, reset_i,
                   output logic sel_i, sel_o, sel_b, rd_addr, wr_addr, enables, read_o, write_o, reset_o
                   );
                   
                   // WIRES
                   logic count_increase;
                   logic result;
                   logic rst;
                   
                   ControlFSM FSM (.clk, .result, .rst, .we(enables), .incr(count_increase));
                   
                   counter COUNT (.clk, .rst, .enb(count_increase), .q(rd_addr));
endmodule
